/****************************************************************************************

	File name    : 
	LastEditors  : H
	LastEditTime : 2021-09-26 18:24:40
	Last Version : 1.0
	Description  : 
	
	----------------------------------------------------------------------------------------
	
	Author       : H
	Date         : 2021-09-26 18:24:39
	FilePath     : \MIPS_32_bit\half_adder.v
	Copyright 2021 H, All Rights Reserved. 

****************************************************************************************/
`ifndef _half_adder
`define _half_adder

module half_adder (
    input   a,
    input   b
    
);
    
endmodule

`endif 