/****************************************************************************************

	File name    : CLA_32_bits_adder
	LastEditors  : H
	LastEditTime : 2021-09-26 19:50:39
	Last Version : 1.0
	Description  : 
	
	----------------------------------------------------------------------------------------
	
	Author       : H
	Date         : 2021-09-26 19:50:37
	FilePath     : \MIPS_32_bit\CLA_adder\CLA_32_bits_adder.v
	Copyright 2021 H, All Rights Reserved. 

****************************************************************************************/
module CLA_32_bits_adder (
    input   [31:0]      A,
    input   [31:0]      B,
    input               Cin,
    
    output              Cout,
    output  [31:0]      S
);
    
endmodule