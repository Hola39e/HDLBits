/****************************************************************************************

	File name    : Control_Unit.v
	LastEditors  : H
	LastEditTime : 2021-09-25 12:21:26
	Last Version : 1.0
	Description  : 
	
	----------------------------------------------------------------------------------------
	
	Author       : H
	Date         : 2021-09-25 12:21:24
	FilePath     : \RISCV_Project\rtl\Control_Unit.v
	Copyright 2021 H, All Rights Reserved. 

****************************************************************************************/
module Control_Unit (
    input   [3:0]   opcode,
    output  reg [1:0]   alu_op,
    output  reg         jump,
                        beq,
                        bne,
                        mem_read,
                        mem_write,
                        alu_src,
                        reg_dst,
                        mem_to_reg,
                        reg_write
);
    always @(*) begin
        case (opcode)
            4'b0000: begin
                reg_dst = 1'b0;
                alu_src = 1'b1;
                mem_to_reg = 1'b1;
                reg_write = 1'b1;
                mem_read = 1'b1;
                mem_write = 1'b0;
                beq = 1'b0;
                bne = 1'b0;
                alu_op = 2'b10;
                jump = 1'b0;   
            end
             4'b0001:  // SW
                begin
                    reg_dst = 1'b0;
                    alu_src = 1'b1;
                    mem_to_reg = 1'b0;
                    reg_write = 1'b0;
                    mem_read = 1'b0;
                    mem_write = 1'b1;
                    beq = 1'b0;
                    bne = 1'b0;
                    alu_op = 2'b10;
                    jump = 1'b0;   
                end
            4'b0010:  // data_processing
                begin
                    reg_dst = 1'b1;
                    alu_src = 1'b0;
                    mem_to_reg = 1'b0;
                    reg_write = 1'b1;
                    mem_read = 1'b0;
                    mem_write = 1'b0;
                    beq = 1'b0;
                    bne = 1'b0;
                    alu_op = 2'b00;
                    jump = 1'b0;   
                end
            4'b0011:  // data_processing
                begin
                    reg_dst = 1'b1;
                    alu_src = 1'b0;
                    mem_to_reg = 1'b0;
                    reg_write = 1'b1;
                    mem_read = 1'b0;
                    mem_write = 1'b0;
                    beq = 1'b0;
                    bne = 1'b0;
                    alu_op = 2'b00;
                    jump = 1'b0;   
                end
            4'b0100:  // data_processing
                begin
                    reg_dst = 1'b1;
                    alu_src = 1'b0;
                    mem_to_reg = 1'b0;
                    reg_write = 1'b1;
                    mem_read = 1'b0;
                    mem_write = 1'b0;
                    beq = 1'b0;
                    bne = 1'b0;
                    alu_op = 2'b00;
                    jump = 1'b0;   
                end
            4'b0101:  // data_processing
                begin
                    reg_dst = 1'b1;
                    alu_src = 1'b0;
                    mem_to_reg = 1'b0;
                    reg_write = 1'b1;
                    mem_read = 1'b0;
                    mem_write = 1'b0;
                    beq = 1'b0;
                    bne = 1'b0;
                    alu_op = 2'b00;
                    jump = 1'b0;   
                end
            4'b0101:  // data_processing
                begin
                    reg_dst = 1'b1;
                    alu_src = 1'b0;
                    mem_to_reg = 1'b0;
                    reg_write = 1'b1;
                    mem_read = 1'b0;
                    mem_write = 1'b0;
                    beq = 1'b0;
                    bne = 1'b0;
                    alu_op = 2'b00;
                    jump = 1'b0;   
                end
            4'b0110:  // data_processing
                begin
                    reg_dst = 1'b1;
                    alu_src = 1'b0;
                    mem_to_reg = 1'b0;
                    reg_write = 1'b1;
                    mem_read = 1'b0;
                    mem_write = 1'b0;
                    beq = 1'b0;
                    bne = 1'b0;
                    alu_op = 2'b00;
                    jump = 1'b0;   
                end
            4'b0111:  // data_processing
                begin
                    reg_dst = 1'b1;
                    alu_src = 1'b0;
                    mem_to_reg = 1'b0;
                    reg_write = 1'b1;
                    mem_read = 1'b0;
                    mem_write = 1'b0;
                    beq = 1'b0;
                    bne = 1'b0;
                    alu_op = 2'b00;
                    jump = 1'b0;   
                end
            4'b1000:  // data_processing
                begin
                    reg_dst = 1'b1;
                    alu_src = 1'b0;
                    mem_to_reg = 1'b0;
                    reg_write = 1'b1;
                    mem_read = 1'b0;
                    mem_write = 1'b0;
                    beq = 1'b0;
                    bne = 1'b0;
                    alu_op = 2'b00;
                    jump = 1'b0;   
                end
            4'b1001:  // data_processing
                begin
                    reg_dst = 1'b1;
                    alu_src = 1'b0;
                    mem_to_reg = 1'b0;
                    reg_write = 1'b1;
                    mem_read = 1'b0;
                    mem_write = 1'b0;
                    beq = 1'b0;
                    bne = 1'b0;
                    alu_op = 2'b00;
                    jump = 1'b0;   
                end
            4'b1011:  // BEQ
                begin
                    reg_dst = 1'b0;
                    alu_src = 1'b0;
                    mem_to_reg = 1'b0;
                    reg_write = 1'b0;
                    mem_read = 1'b0;
                    mem_write = 1'b0;
                    beq = 1'b1;
                    bne = 1'b0;
                    alu_op = 2'b01;
                    jump = 1'b0;   
                end
            4'b1100:  // BNE
                begin
                    reg_dst = 1'b0;
                    alu_src = 1'b0;
                    mem_to_reg = 1'b0;
                    reg_write = 1'b0;
                    mem_read = 1'b0;
                    mem_write = 1'b0;
                    beq = 1'b0;
                    bne = 1'b1;
                    alu_op = 2'b01;
                    jump = 1'b0;   
                end
            4'b1101:  // J
                begin
                    reg_dst = 1'b0;
                    alu_src = 1'b0;
                    mem_to_reg = 1'b0;
                    reg_write = 1'b0;
                    mem_read = 1'b0;
                    mem_write = 1'b0;
                    beq = 1'b0;
                    bne = 1'b0;
                    alu_op = 2'b00;
                    jump = 1'b1;   
                end   
            default: begin
                    reg_dst = 1'b1;
                    alu_src = 1'b0;
                    mem_to_reg = 1'b0;
                    reg_write = 1'b1;
                    mem_read = 1'b0;
                    mem_write = 1'b0;
                    beq = 1'b0;
                    bne = 1'b0;
                    alu_op = 2'b00;
                    jump = 1'b0; 
                end
        endcase
    end
endmodule